module bitwise_invert(a, out);
input [31:0] a;
output [31:0] out;

not not0(out[0], a[0]);
not not1(out[1], a[1]);
not not2(out[2], a[2]);
not not3(out[3], a[3]);
not not4(out[4], a[4]);
not not5(out[5], a[5]);
not not6(out[6], a[6]);
not not7(out[7], a[7]);
not not8(out[8], a[8]);
not not9(out[9], a[9]);
not not10(out[10], a[10]);
not not11(out[11], a[11]);
not not12(out[12], a[12]);
not not13(out[13], a[13]);
not not14(out[14], a[14]);
not not15(out[15], a[15]);
not not16(out[16], a[16]);
not not17(out[17], a[17]);
not not18(out[18], a[18]);
not not19(out[19], a[19]);
not not20(out[20], a[20]);
not not21(out[21], a[21]);
not not22(out[22], a[22]);
not not23(out[23], a[23]);
not not24(out[24], a[24]);
not not25(out[25], a[25]);
not not26(out[26], a[26]);
not not27(out[27], a[27]);
not not28(out[28], a[28]);
not not29(out[29], a[29]);
not not30(out[30], a[30]);
not not31(out[31], a[31]);
endmodule